/*
 * Copyright (c) 2011-2012 Travis Geiselbrecht
 *
 * Permission is hereby granted, free of charge, to any person obtaining
 * a copy of this software and associated documentation files
 * (the "Software"), to deal in the Software without restriction,
 * including without limitation the rights to use, copy, modify, merge,
 * publish, distribute, sublicense, and/or sell copies of the Software,
 * and to permit persons to whom the Software is furnished to do so,
 * subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be
 * included in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
 * EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
 * MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
 * IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
 * CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
 * TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
 * SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 */
module top
	(
		////////////////////	Clock Input	 	////////////////////	 
		CLOCK_24,						//	24 MHz
		CLOCK_27,						//	27 MHz
		CLOCK_50,						//	50 MHz
		EXT_CLOCK,						//	External Clock
		////////////////////	Push Button		////////////////////
		KEY,							//	Pushbutton[3:0]
		////////////////////	DPDT Switch		////////////////////
		SW,								//	Toggle Switch[9:0]
		////////////////////	7-SEG Dispaly	////////////////////
		HEX0,							//	Seven Segment Digit 0
		HEX1,							//	Seven Segment Digit 1
		HEX2,							//	Seven Segment Digit 2
		HEX3,							//	Seven Segment Digit 3
		////////////////////////	LED		////////////////////////
		LEDG,							//	LED Green[7:0]
		LEDR,							//	LED Red[9:0]
		////////////////////////	UART	////////////////////////
		UART_TXD,						//	UART Transmitter
		UART_RXD,						//	UART Receiver
		/////////////////////	SDRAM Interface		////////////////
		DRAM_DQ,						//	SDRAM Data bus 16 Bits
		DRAM_ADDR,						//	SDRAM Address bus 12 Bits
		DRAM_LDQM,						//	SDRAM Low-byte Data Mask 
		DRAM_UDQM,						//	SDRAM High-byte Data Mask
		DRAM_WE_N,						//	SDRAM Write Enable
		DRAM_CAS_N,						//	SDRAM Column Address Strobe
		DRAM_RAS_N,						//	SDRAM Row Address Strobe
		DRAM_CS_N,						//	SDRAM Chip Select
		DRAM_BA_0,						//	SDRAM Bank Address 0
		DRAM_BA_1,						//	SDRAM Bank Address 0
		DRAM_CLK,						//	SDRAM Clock
		DRAM_CKE,						//	SDRAM Clock Enable
		////////////////////	Flash Interface		////////////////
		FL_DQ,							//	FLASH Data bus 8 Bits
		FL_ADDR,						//	FLASH Address bus 22 Bits
		FL_WE_N,						//	FLASH Write Enable
		FL_RST_N,						//	FLASH Reset
		FL_OE_N,						//	FLASH Output Enable
		FL_CE_N,						//	FLASH Chip Enable
		////////////////////	SRAM Interface		////////////////
		SRAM_DQ,						//	SRAM Data bus 16 Bits
		SRAM_ADDR,						//	SRAM Address bus 18 Bits
		SRAM_UB_N,						//	SRAM High-byte Data Mask 
		SRAM_LB_N,						//	SRAM Low-byte Data Mask 
		SRAM_WE_N,						//	SRAM Write Enable
		SRAM_CE_N,						//	SRAM Chip Enable
		SRAM_OE_N,						//	SRAM Output Enable
		////////////////////	SD_Card Interface	////////////////
		SD_DAT,							//	SD Card Data
		SD_DAT3,						//	SD Card Data 3
		SD_CMD,							//	SD Card Command Signal
		SD_CLK,							//	SD Card Clock
		////////////////////	USB JTAG link	////////////////////
		TDI,  							// CPLD -> FPGA (data in)
		TCK,  							// CPLD -> FPGA (clk)
		TCS,  							// CPLD -> FPGA (CS)
	    TDO,  							// FPGA -> CPLD (data out)
		////////////////////	I2C		////////////////////////////
		I2C_SDAT,						//	I2C Data
		I2C_SCLK,						//	I2C Clock
		////////////////////	PS2		////////////////////////////
		PS2_DAT,						//	PS2 Data
		PS2_CLK,						//	PS2 Clock
		////////////////////	VGA		////////////////////////////
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_R,   						//	VGA Red[3:0]
		VGA_G,	 						//	VGA Green[3:0]
		VGA_B,  						//	VGA Blue[3:0]
		////////////////	Audio CODEC		////////////////////////
		AUD_ADCLRCK,					//	Audio CODEC ADC LR Clock
		AUD_ADCDAT,						//	Audio CODEC ADC Data
		AUD_DACLRCK,					//	Audio CODEC DAC LR Clock
		AUD_DACDAT,						//	Audio CODEC DAC Data
		AUD_BCLK,						//	Audio CODEC Bit-Stream Clock
		AUD_XCK,						//	Audio CODEC Chip Clock
		////////////////////	GPIO	////////////////////////////
		GPIO_0,							//	GPIO Connection 0
		GPIO_1							//	GPIO Connection 1
	);

////////////////////////	Clock Input	 	////////////////////////
input	[1:0]	CLOCK_24;				//	24 MHz
input	[1:0]	CLOCK_27;				//	27 MHz
input			CLOCK_50;				//	50 MHz
input			EXT_CLOCK;				//	External Clock
////////////////////////	Push Button		////////////////////////
input	[3:0]	KEY;					//	Pushbutton[3:0]
////////////////////////	DPDT Switch		////////////////////////
input	[9:0]	SW;						//	Toggle Switch[9:0]
////////////////////////	7-SEG Dispaly	////////////////////////
output	[6:0]	HEX0;					//	Seven Segment Digit 0
output	[6:0]	HEX1;					//	Seven Segment Digit 1
output	[6:0]	HEX2;					//	Seven Segment Digit 2
output	[6:0]	HEX3;					//	Seven Segment Digit 3
////////////////////////////	LED		////////////////////////////
output	[7:0]	LEDG;					//	LED Green[7:0]
output	[9:0]	LEDR;					//	LED Red[9:0]
////////////////////////////	UART	////////////////////////////
output			UART_TXD;				//	UART Transmitter
input			UART_RXD;				//	UART Receiver
///////////////////////		SDRAM Interface	////////////////////////
inout	[15:0]	DRAM_DQ;				//	SDRAM Data bus 16 Bits
output	[11:0]	DRAM_ADDR;				//	SDRAM Address bus 12 Bits
output			DRAM_LDQM;				//	SDRAM Low-byte Data Mask 
output			DRAM_UDQM;				//	SDRAM High-byte Data Mask
output			DRAM_WE_N;				//	SDRAM Write Enable
output			DRAM_CAS_N;				//	SDRAM Column Address Strobe
output			DRAM_RAS_N;				//	SDRAM Row Address Strobe
output			DRAM_CS_N;				//	SDRAM Chip Select
output			DRAM_BA_0;				//	SDRAM Bank Address 0
output			DRAM_BA_1;				//	SDRAM Bank Address 0
output			DRAM_CLK;				//	SDRAM Clock
output			DRAM_CKE;				//	SDRAM Clock Enable
////////////////////////	Flash Interface	////////////////////////
inout	[7:0]	FL_DQ;					//	FLASH Data bus 8 Bits
output	[21:0]	FL_ADDR;				//	FLASH Address bus 22 Bits
output			FL_WE_N;				//	FLASH Write Enable
output			FL_RST_N;				//	FLASH Reset
output			FL_OE_N;				//	FLASH Output Enable
output			FL_CE_N;				//	FLASH Chip Enable
////////////////////////	SRAM Interface	////////////////////////
inout	[15:0]	SRAM_DQ;				//	SRAM Data bus 16 Bits
output	[17:0]	SRAM_ADDR;				//	SRAM Address bus 18 Bits
output			SRAM_UB_N;				//	SRAM High-byte Data Mask 
output			SRAM_LB_N;				//	SRAM Low-byte Data Mask 
output			SRAM_WE_N;				//	SRAM Write Enable
output			SRAM_CE_N;				//	SRAM Chip Enable
output			SRAM_OE_N;				//	SRAM Output Enable
////////////////////	SD Card Interface	////////////////////////
inout			SD_DAT;					//	SD Card Data
inout			SD_DAT3;				//	SD Card Data 3
inout			SD_CMD;					//	SD Card Command Signal
output			SD_CLK;					//	SD Card Clock
////////////////////////	I2C		////////////////////////////////
inout			I2C_SDAT;				//	I2C Data
output			I2C_SCLK;				//	I2C Clock
////////////////////////	PS2		////////////////////////////////
input		 	PS2_DAT;				//	PS2 Data
input			PS2_CLK;				//	PS2 Clock
////////////////////	USB JTAG link	////////////////////////////
input  			TDI;					// CPLD -> FPGA (data in)
input  			TCK;					// CPLD -> FPGA (clk)
input  			TCS;					// CPLD -> FPGA (CS)
output 			TDO;					// FPGA -> CPLD (data out)
////////////////////////	VGA			////////////////////////////
output			VGA_HS;					//	VGA H_SYNC
output			VGA_VS;					//	VGA V_SYNC
output	[3:0]	VGA_R;   				//	VGA Red[3:0]
output	[3:0]	VGA_G;	 				//	VGA Green[3:0]
output	[3:0]	VGA_B;   				//	VGA Blue[3:0]
////////////////////	Audio CODEC		////////////////////////////
output			AUD_ADCLRCK;			//	Audio CODEC ADC LR Clock
input			AUD_ADCDAT;				//	Audio CODEC ADC Data
output			AUD_DACLRCK;			//	Audio CODEC DAC LR Clock
output			AUD_DACDAT;				//	Audio CODEC DAC Data
inout			AUD_BCLK;				//	Audio CODEC Bit-Stream Clock
output			AUD_XCK;				//	Audio CODEC Chip Clock
////////////////////////	GPIO	////////////////////////////////
input	[35:0]	GPIO_0;					//	GPIO Connection 0
inout	[35:0]	GPIO_1;					//	GPIO Connection 1
///////////////////////////////////////////////////////////////////

//assign GPIO_1 = GPIO_0;

// run a 1mhz clock
reg[6:0] div;

initial begin
	div <= 0;
end

always @(posedge CLOCK_24[0])
begin
	div = div + 1;
end

wire slowclk = CLOCK_24[0]; //div[4];

/*
reg slowclk;
always @(negedge KEY[0])
begin
	slowclk <= ~slowclk;
end
*/

/* instantiate the cpu */
wire cpu_re;
wire cpu_we;
reg rst;
wire [29:0] memaddr;
wire [31:0] rmemdata;
wire [31:0] wmemdata;
wire [31:0] cpudebugout;

//assign rst = KEY[0];

initial
	rst <= 0;

cpu cpu0(
	.clk(slowclk),
	.rst(rst),
	.mem_re(cpu_re),
	.mem_we(cpu_we),
	.memaddr(memaddr),
	.rmemdata(rmemdata),
	.wmemdata(wmemdata),

	.debugout(cpudebugout)
);

/* main memory */
wire mem_re = cpu_re && (memaddr[29] == 0);
wire mem_we = cpu_we && (memaddr[29] == 0);

syncmem mem0(
	.clk(slowclk),
	.re(mem_re),
	.we(mem_we),
	.addr(memaddr),
	.rdata(rmemdata),
	.wdata(wmemdata)
);

/* uart */
wire uart_re = cpu_re && (memaddr[29:14] == 16'b1000000000000000);
wire uart_we = cpu_we && (memaddr[29:14] == 16'b1000000000000000);

uart uart0(
	.clk(slowclk),
	.rst(rst),

	.hwtx(UART_TXD),
	.hwrx(UART_RXD),

	.addr(memaddr[0]),
	.re(uart_re),
	.we(uart_we),
	.wdata(wmemdata),
	.rdata(rmemdata),

//	.rxchar(0),
//	.rxvalid(),
	);

/* debug register */
wire debuglatch_we = cpu_we && (memaddr[29:14] == 16'b1000000000000001);

reg[31:0] debuglatch;
always @(posedge slowclk) begin
	if (debuglatch_we) begin
		debuglatch <= wmemdata;
	end
end


//`define WITH_SRAM
`ifdef WITH_SRAM
assign SRAM_UB_N = 0;
assign SRAM_LB_N = 0;

wire read_sync;
wire write_sync;

integer addr;

reg [1:0] retest;
always @(negedge slowclk) begin
	retest <= retest + 1;
end

always @(posedge read_sync or posedge write_sync) begin
	addr <= addr + 1;
end

sramcontroller sram(
	.clk(slowclk),
	.addr(addr),
	.indata(0),
	.re(retest[1]),
	.we(retest[0]),
	.read_sync(read_sync),
	.write_sync(write_sync),

	.memclk(memclk),
	.sram_addr(SRAM_ADDR),
	.sram_data(SRAM_DQ),
	.sram_ce(SRAM_CE_N),
	.sram_re(SRAM_OE_N),
	.sram_we(SRAM_WE_N)
);
`endif

reg[15:0] debugreg;

always @(SW[9] or SW[8] or SW[7] or memaddr or rmemdata or debuglatch)
begin
	if (SW[9]) begin
		debugreg = rmemdata[31:16];
	end else if (SW[8]) begin
		debugreg = rmemdata[15:0];
	end else if (SW[7]) begin
		debugreg = memaddr[29:16];
	end else if (SW[1]) begin
		debugreg = debuglatch[31:16];
	end else if (SW[0]) begin
		debugreg = debuglatch[15:0];
	end else begin
		debugreg = memaddr[15:0];
	end
end

/* debug info */
seven_segment seg0(debugreg[3:0], HEX0);
seven_segment seg1(debugreg[7:4], HEX1);
seven_segment seg2(debugreg[11:8], HEX2);
seven_segment seg3(debugreg[15:12], HEX3);

assign LEDG[0] = rst;
assign LEDG[1] = slowclk;
assign LEDG[2] = mem_re;
assign LEDG[3] = mem_we;

//assign GPIO_1[0] = slowclk;
//assign GPIO_1[1] = mem_re;
//assign GPIO_1[2] = mem_we;
//assign GPIO_1[7:3] = memaddr[4:0];

//assign GPIO_1[15:8] = wmemdata[7:0];
//assign GPIO_1[8] = memclk;
//assign GPIO_1[9] = read_sync;
//assign GPIO_1[10] = write_sync;
//assign GPIO_1[11] = SRAM_CE_N;
//assign GPIO_1[12] = SRAM_OE_N;
//assign GPIO_1[15:13] = SRAM_ADDR[2:0];

assign GPIO_1[0] = UART_TXD;
assign GPIO_1[1] = UART_RXD;

endmodule

module syncmem(
	input clk,
	input re,
	input we,
	input [29:0] addr,
	output reg [31:0] rdata,
	input [31:0] wdata
);

reg [31:0] mem [0:4096];

initial begin
	$readmemh("../test/test2.asm.hex", mem);
end

always @(posedge clk) begin
	if (re)
		rdata <= mem[addr];
	else
		rdata <= 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
	if (we)
		mem[addr] <= wdata;
end

endmodule

